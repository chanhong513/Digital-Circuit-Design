module convolution_3by3_module (
    // Inputs
    clk,
    rst,
    buffer_read_addr_in_3by3,
    input_side_array_addr_in_3by3, input_ceiling_array_addr_in_3by3, filter_side_array_addr_in_3by3, filter_ceiling_array_addr_in_3by3,
    sys_3by3_en,

    a00_output, a01_output, a02_output, a03_output, 
    a10_output, a11_output, a12_output, a13_output, 
    a20_output, a21_output, a22_output, a23_output, 
    a30_output, a31_output, a32_output, a33_output, 
    b00_output, b01_output, b02_output, 
    b10_output, b11_output, b12_output, 
    b20_output, b21_output, b22_output, 
    zero_input,
    

    // Outputs
    convolution_C11,
    convolution_C12,
    convolution_C21,
    convolution_C22,

    convolution_3by3_out
    );

    // input
    input clk;
    input rst;
    input [1:0] buffer_read_addr_in_3by3;
    input [4:0] input_side_array_addr_in_3by3, input_ceiling_array_addr_in_3by3, filter_side_array_addr_in_3by3, filter_ceiling_array_addr_in_3by3;
    input sys_3by3_en;
    input [7:0] a00_output, a01_output, a02_output, a03_output, a10_output, a11_output, a12_output, a13_output, a20_output, a21_output, a22_output, a23_output, a30_output, a31_output, a32_output, a33_output, b00_output, b01_output, b02_output, b10_output, b11_output, b12_output, b20_output, b21_output, b22_output, zero_input;
    
    // output wire [4:0] state_output, next_state_output;
    output wire [7:0] convolution_3by3_out;
    output wire [7:0] convolution_C11, convolution_C12, convolution_C21, convolution_C22;


    // Instantiate the MUX
    wire [7:0] out_side_input;
    // output wire [4:0] sel_input;
    MUX_32bit mux_3by3_input_side (
        .i0(a00_output), .i1(a01_output), .i2(a02_output), .i3(a03_output), .i4(a10_output), .i5(a11_output), .i6(a12_output), .i7(a13_output),
        .i8(a20_output), .i9(a21_output), .i10(a22_output), .i11(a23_output), .i12(a30_output), .i13(a31_output), .i14(a32_output), .i15(a33_output),
        .i16(b00_output), .i17(b01_output), .i18(b02_output), .i19(b10_output), .i20(b11_output), .i21(b12_output), .i22(b20_output), .i23(b21_output), .i24(b22_output), 
        .i25(zero_input), .i26(8'b0), .i27(8'b0), .i28(8'b0), .i29(8'b0), .i30(8'b0), .i31(8'b0),
        .sel(input_side_array_addr_in_3by3),
        .out(out_side_input)
    );

    // Instantiate the MUX
    wire [7:0] out_ceiling_input;
    // output wire [4:0] sel_input;
    MUX_32bit mux_3by3_input_ceiling (
        .i0(a00_output), .i1(a01_output), .i2(a02_output), .i3(a03_output), .i4(a10_output), .i5(a11_output), .i6(a12_output), .i7(a13_output),
        .i8(a20_output), .i9(a21_output), .i10(a22_output), .i11(a23_output), .i12(a30_output), .i13(a31_output), .i14(a32_output), .i15(a33_output),
        .i16(b00_output), .i17(b01_output), .i18(b02_output), .i19(b10_output), .i20(b11_output), .i21(b12_output), .i22(b20_output), .i23(b21_output), .i24(b22_output), 
        .i25(zero_input), .i26(8'b0), .i27(8'b0), .i28(8'b0), .i29(8'b0), .i30(8'b0), .i31(8'b0),
        .sel(input_ceiling_array_addr_in_3by3),
        .out(out_ceiling_input)
    );

    // Instantiate the MUX
    wire [7:0] out_side_filter;
    // output wire [4:0] filter_side_array_addr_in_3by3;
    MUX_32bit mux_3by3_side_filter (
        .i0(a00_output), .i1(a01_output), .i2(a02_output), .i3(a03_output), .i4(a10_output), .i5(a11_output), .i6(a12_output), .i7(a13_output),
        .i8(a20_output), .i9(a21_output), .i10(a22_output), .i11(a23_output), .i12(a30_output), .i13(a31_output), .i14(a32_output), .i15(a33_output),
        .i16(b00_output), .i17(b01_output), .i18(b02_output), .i19(b10_output), .i20(b11_output), .i21(b12_output), .i22(b20_output), .i23(b21_output), .i24(b22_output), 
        .i25(zero_input), .i26(8'b0), .i27(8'b0), .i28(8'b0), .i29(8'b0), .i30(8'b0), .i31(8'b0),
        .sel(filter_side_array_addr_in_3by3),
        .out(out_side_filter)
    );

    // Instantiate the MUX
    wire [7:0] out_ceiling_filter;
    // output wire [4:0] filter_ceiling_array_addr_in_3by3;
    MUX_32bit mux_3by3_ceiling_filter (
        .i0(a00_output), .i1(a01_output), .i2(a02_output), .i3(a03_output), .i4(a10_output), .i5(a11_output), .i6(a12_output), .i7(a13_output),
        .i8(a20_output), .i9(a21_output), .i10(a22_output), .i11(a23_output), .i12(a30_output), .i13(a31_output), .i14(a32_output), .i15(a33_output),
        .i16(b00_output), .i17(b01_output), .i18(b02_output), .i19(b10_output), .i20(b11_output), .i21(b12_output), .i22(b20_output), .i23(b21_output), .i24(b22_output), 
        .i25(zero_input), .i26(8'b0), .i27(8'b0), .i28(8'b0), .i29(8'b0), .i30(8'b0), .i31(8'b0),
        .sel(filter_ceiling_array_addr_in_3by3),
        .out(out_ceiling_filter)
    );


    // output wire [7:0] side_1, side_2, ceiling_1, ceiling_2;
    // Instantiate the Systolic_Array_2x2_module
    Systolic_Array_3x3_module systolic_array_3x3 (
        .clk(clk), 
        .rst(rst),
        .en(sys_3by3_en),
        .side_1(out_side_input),
        .side_2(out_side_input),
        .side_3(out_side_filter),
        .ceiling_1(out_ceiling_filter),
        .ceiling_2(out_ceiling_input),
        .ceiling_3(out_ceiling_input),
        .convolution_11(convolution_C11),
        .convolution_12(convolution_C12),
        .convolution_21(convolution_C21),
        .convolution_22(convolution_C22)
    );


    buffer_module buffer_3by3(
        .clk(clk),
        .rst(rst),
        .buffer_read_addr_in(buffer_read_addr_in_3by3), // 2bits
        .data_in_0(convolution_C11), // 8bits
        .data_in_1(convolution_C12), // 8bits
        .data_in_2(convolution_C21), // 8bits
        .data_in_3(convolution_C22), // 8bits
        .data_out(convolution_3by3_out) // 8bits
    );

endmodule
